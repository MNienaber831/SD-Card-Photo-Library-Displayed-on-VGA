// nios_system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module nios_system (
		input  wire [3:0]  pushbuttons_export,         //          pushbuttons.export
		inout  wire        sd_card_b_SD_cmd,           //              sd_card.b_SD_cmd
		inout  wire        sd_card_b_SD_dat,           //                     .b_SD_dat
		inout  wire        sd_card_b_SD_dat3,          //                     .b_SD_dat3
		output wire        sd_card_o_SD_clock,         //                     .o_SD_clock
		output wire [12:0] sdram_addr,                 //                sdram.addr
		output wire [1:0]  sdram_ba,                   //                     .ba
		output wire        sdram_cas_n,                //                     .cas_n
		output wire        sdram_cke,                  //                     .cke
		output wire        sdram_cs_n,                 //                     .cs_n
		inout  wire [15:0] sdram_dq,                   //                     .dq
		output wire [1:0]  sdram_dqm,                  //                     .dqm
		output wire        sdram_ras_n,                //                     .ras_n
		output wire        sdram_we_n,                 //                     .we_n
		output wire        sdram_clk_clk,              //            sdram_clk.clk
		inout  wire [15:0] sram_DQ,                    //                 sram.DQ
		output wire [19:0] sram_ADDR,                  //                     .ADDR
		output wire        sram_LB_N,                  //                     .LB_N
		output wire        sram_UB_N,                  //                     .UB_N
		output wire        sram_CE_N,                  //                     .CE_N
		output wire        sram_OE_N,                  //                     .OE_N
		output wire        sram_WE_N,                  //                     .WE_N
		input  wire        system_pll_ref_clk_clk,     //   system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset, // system_pll_ref_reset.reset
		output wire        vga_CLK,                    //                  vga.CLK
		output wire        vga_HS,                     //                     .HS
		output wire        vga_VS,                     //                     .VS
		output wire        vga_BLANK,                  //                     .BLANK
		output wire        vga_SYNC,                   //                     .SYNC
		output wire [7:0]  vga_R,                      //                     .R
		output wire [7:0]  vga_G,                      //                     .G
		output wire [7:0]  vga_B,                      //                     .B
		input  wire        vga_pll_ref_clk_clk,        //      vga_pll_ref_clk.clk
		input  wire        vga_pll_ref_reset_reset     //    vga_pll_ref_reset.reset
	);

	wire         system_pll_sys_clk_clk;                                             // System_PLL:sys_clk_clk -> [Interval_Timer:clk, JTAG_UART:clk, Nios2:clk, Pushbuttons:clk, SDRAM:clk, SD_Card:i_clock, SRAM:clk, SysID:clock, VGA_Subsystem:sys_clk_clk, irq_mapper:clk, mm_interconnect_0:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_001:clk]
	wire         system_pll_reset_source_reset;                                      // System_PLL:reset_source_reset -> [VGA_Subsystem:sys_reset_reset_n, rst_controller:reset_in0, rst_controller_001:reset_in1]
	wire  [31:0] nios2_data_master_readdata;                                         // mm_interconnect_0:Nios2_data_master_readdata -> Nios2:d_readdata
	wire         nios2_data_master_waitrequest;                                      // mm_interconnect_0:Nios2_data_master_waitrequest -> Nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                      // Nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Nios2_data_master_debugaccess
	wire  [27:0] nios2_data_master_address;                                          // Nios2:d_address -> mm_interconnect_0:Nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                       // Nios2:d_byteenable -> mm_interconnect_0:Nios2_data_master_byteenable
	wire         nios2_data_master_read;                                             // Nios2:d_read -> mm_interconnect_0:Nios2_data_master_read
	wire         nios2_data_master_readdatavalid;                                    // mm_interconnect_0:Nios2_data_master_readdatavalid -> Nios2:d_readdatavalid
	wire         nios2_data_master_write;                                            // Nios2:d_write -> mm_interconnect_0:Nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                        // Nios2:d_writedata -> mm_interconnect_0:Nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                                  // mm_interconnect_0:Nios2_instruction_master_readdata -> Nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                               // mm_interconnect_0:Nios2_instruction_master_waitrequest -> Nios2:i_waitrequest
	wire  [27:0] nios2_instruction_master_address;                                   // Nios2:i_address -> mm_interconnect_0:Nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                      // Nios2:i_read -> mm_interconnect_0:Nios2_instruction_master_read
	wire         nios2_instruction_master_readdatavalid;                             // mm_interconnect_0:Nios2_instruction_master_readdatavalid -> Nios2:i_readdatavalid
	wire         vga_subsystem_pixel_dma_master_waitrequest;                         // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_waitrequest -> VGA_Subsystem:pixel_dma_master_waitrequest
	wire  [15:0] vga_subsystem_pixel_dma_master_readdata;                            // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdata -> VGA_Subsystem:pixel_dma_master_readdata
	wire  [31:0] vga_subsystem_pixel_dma_master_address;                             // VGA_Subsystem:pixel_dma_master_address -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_address
	wire         vga_subsystem_pixel_dma_master_read;                                // VGA_Subsystem:pixel_dma_master_read -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_read
	wire         vga_subsystem_pixel_dma_master_readdatavalid;                       // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdatavalid -> VGA_Subsystem:pixel_dma_master_readdatavalid
	wire         vga_subsystem_pixel_dma_master_lock;                                // VGA_Subsystem:pixel_dma_master_lock -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_lock
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;           // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;             // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;          // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;              // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                 // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;            // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect;           // mm_interconnect_0:SD_Card_avalon_sdcard_slave_chipselect -> SD_Card:i_avalon_chip_select
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata;             // SD_Card:o_avalon_readdata -> mm_interconnect_0:SD_Card_avalon_sdcard_slave_readdata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest;          // SD_Card:o_avalon_waitrequest -> mm_interconnect_0:SD_Card_avalon_sdcard_slave_waitrequest
	wire   [7:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_address;              // mm_interconnect_0:SD_Card_avalon_sdcard_slave_address -> SD_Card:i_avalon_address
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_read;                 // mm_interconnect_0:SD_Card_avalon_sdcard_slave_read -> SD_Card:i_avalon_read
	wire   [3:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable;           // mm_interconnect_0:SD_Card_avalon_sdcard_slave_byteenable -> SD_Card:i_avalon_byteenable
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_write;                // mm_interconnect_0:SD_Card_avalon_sdcard_slave_write -> SD_Card:i_avalon_write
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata;            // mm_interconnect_0:SD_Card_avalon_sdcard_slave_writedata -> SD_Card:i_avalon_writedata
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_readdata;                  // SRAM:readdata -> mm_interconnect_0:SRAM_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_sram_slave_address;                   // mm_interconnect_0:SRAM_avalon_sram_slave_address -> SRAM:address
	wire         mm_interconnect_0_sram_avalon_sram_slave_read;                      // mm_interconnect_0:SRAM_avalon_sram_slave_read -> SRAM:read
	wire   [1:0] mm_interconnect_0_sram_avalon_sram_slave_byteenable;                // mm_interconnect_0:SRAM_avalon_sram_slave_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_avalon_sram_slave_readdatavalid;             // SRAM:readdatavalid -> mm_interconnect_0:SRAM_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_avalon_sram_slave_write;                     // mm_interconnect_0:SRAM_avalon_sram_slave_write -> SRAM:write
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_writedata;                 // mm_interconnect_0:SRAM_avalon_sram_slave_writedata -> SRAM:writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                     // SysID:readdata -> mm_interconnect_0:SysID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                      // mm_interconnect_0:SysID_control_slave_address -> SysID:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;                   // Nios2:debug_mem_slave_readdata -> mm_interconnect_0:Nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;                // Nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:Nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;                // mm_interconnect_0:Nios2_debug_mem_slave_debugaccess -> Nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;                    // mm_interconnect_0:Nios2_debug_mem_slave_address -> Nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                       // mm_interconnect_0:Nios2_debug_mem_slave_read -> Nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;                 // mm_interconnect_0:Nios2_debug_mem_slave_byteenable -> Nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                      // mm_interconnect_0:Nios2_debug_mem_slave_write -> Nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;                  // mm_interconnect_0:Nios2_debug_mem_slave_writedata -> Nios2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata;   // VGA_Subsystem:pixel_dma_control_slave_readdata -> mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address;    // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_address -> VGA_Subsystem:pixel_dma_control_slave_address
	wire         mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read;       // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_read -> VGA_Subsystem:pixel_dma_control_slave_read
	wire   [3:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable; // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_byteenable -> VGA_Subsystem:pixel_dma_control_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write;      // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_write -> VGA_Subsystem:pixel_dma_control_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata;  // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_writedata -> VGA_Subsystem:pixel_dma_control_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                              // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                             // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                 // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                    // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                              // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                           // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                   // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                               // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_pushbuttons_s1_chipselect;                        // mm_interconnect_0:Pushbuttons_s1_chipselect -> Pushbuttons:chipselect
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_readdata;                          // Pushbuttons:readdata -> mm_interconnect_0:Pushbuttons_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuttons_s1_address;                           // mm_interconnect_0:Pushbuttons_s1_address -> Pushbuttons:address
	wire         mm_interconnect_0_pushbuttons_s1_write;                             // mm_interconnect_0:Pushbuttons_s1_write -> Pushbuttons:write_n
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_writedata;                         // mm_interconnect_0:Pushbuttons_s1_writedata -> Pushbuttons:writedata
	wire         mm_interconnect_0_interval_timer_s1_chipselect;                     // mm_interconnect_0:Interval_Timer_s1_chipselect -> Interval_Timer:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_s1_readdata;                       // Interval_Timer:readdata -> mm_interconnect_0:Interval_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_s1_address;                        // mm_interconnect_0:Interval_Timer_s1_address -> Interval_Timer:address
	wire         mm_interconnect_0_interval_timer_s1_write;                          // mm_interconnect_0:Interval_Timer_s1_write -> Interval_Timer:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_s1_writedata;                      // mm_interconnect_0:Interval_Timer_s1_writedata -> Interval_Timer:writedata
	wire         irq_mapper_receiver0_irq;                                           // Pushbuttons:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                           // Interval_Timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                           // JTAG_UART:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_irq_irq;                                                      // irq_mapper:sender_irq -> Nios2:irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [Interval_Timer:reset_n, JTAG_UART:rst_n, Pushbuttons:reset_n, SDRAM:reset_n, SD_Card:i_reset_n, SRAM:reset, SysID:reset_n, mm_interconnect_0:JTAG_UART_reset_reset_bridge_in_reset_reset, mm_interconnect_0:VGA_Subsystem_sys_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [Nios2:reset_n, irq_mapper:reset, mm_interconnect_0:Nios2_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                             // rst_controller_001:reset_req -> [Nios2:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                                    // Nios2:debug_reset_request -> rst_controller_001:reset_in0

	nios_system_Interval_Timer interval_timer (
		.clk        (system_pll_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                        //   irq.irq
	);

	nios_system_JTAG_UART jtag_uart (
		.clk            (system_pll_sys_clk_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	nios_system_Nios2 nios2 (
		.clk                                 (system_pll_sys_clk_clk),                              //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	nios_system_Pushbuttons pushbuttons (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pushbuttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pushbuttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pushbuttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pushbuttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pushbuttons_s1_readdata),   //                    .readdata
		.in_port    (pushbuttons_export),                          // external_connection.export
		.irq        (irq_mapper_receiver0_irq)                     //                 irq.irq
	);

	nios_system_SDRAM sdram (
		.clk            (system_pll_sys_clk_clk),                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card (
		.i_avalon_chip_select (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (system_pll_sys_clk_clk),                                    //                 clk.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                           //               reset.reset_n
		.b_SD_cmd             (sd_card_b_SD_cmd),                                          //         conduit_end.export
		.b_SD_dat             (sd_card_b_SD_dat),                                          //                    .export
		.b_SD_dat3            (sd_card_b_SD_dat3),                                         //                    .export
		.o_SD_clock           (sd_card_o_SD_clock)                                         //                    .export
	);

	nios_system_SRAM sram (
		.clk           (system_pll_sys_clk_clk),                                 //                clk.clk
		.reset         (rst_controller_reset_out_reset),                         //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                              //                   .export
		.SRAM_LB_N     (sram_LB_N),                                              //                   .export
		.SRAM_UB_N     (sram_UB_N),                                              //                   .export
		.SRAM_CE_N     (sram_CE_N),                                              //                   .export
		.SRAM_OE_N     (sram_OE_N),                                              //                   .export
		.SRAM_WE_N     (sram_WE_N),                                              //                   .export
		.address       (mm_interconnect_0_sram_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	nios_system_SysID sysid (
		.clock    (system_pll_sys_clk_clk),                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	nios_system_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	nios_system_VGA_Subsystem vga_subsystem (
		.pixel_dma_control_slave_address    (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address),    // pixel_dma_control_slave.address
		.pixel_dma_control_slave_byteenable (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable), //                        .byteenable
		.pixel_dma_control_slave_read       (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read),       //                        .read
		.pixel_dma_control_slave_write      (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write),      //                        .write
		.pixel_dma_control_slave_writedata  (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata),  //                        .writedata
		.pixel_dma_control_slave_readdata   (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata),   //                        .readdata
		.pixel_dma_master_readdatavalid     (vga_subsystem_pixel_dma_master_readdatavalid),                       //        pixel_dma_master.readdatavalid
		.pixel_dma_master_waitrequest       (vga_subsystem_pixel_dma_master_waitrequest),                         //                        .waitrequest
		.pixel_dma_master_address           (vga_subsystem_pixel_dma_master_address),                             //                        .address
		.pixel_dma_master_lock              (vga_subsystem_pixel_dma_master_lock),                                //                        .lock
		.pixel_dma_master_read              (vga_subsystem_pixel_dma_master_read),                                //                        .read
		.pixel_dma_master_readdata          (vga_subsystem_pixel_dma_master_readdata),                            //                        .readdata
		.sys_clk_clk                        (system_pll_sys_clk_clk),                                             //                 sys_clk.clk
		.sys_reset_reset_n                  (~system_pll_reset_source_reset),                                     //               sys_reset.reset_n
		.vga_CLK                            (vga_CLK),                                                            //                     vga.CLK
		.vga_HS                             (vga_HS),                                                             //                        .HS
		.vga_VS                             (vga_VS),                                                             //                        .VS
		.vga_BLANK                          (vga_BLANK),                                                          //                        .BLANK
		.vga_SYNC                           (vga_SYNC),                                                           //                        .SYNC
		.vga_R                              (vga_R),                                                              //                        .R
		.vga_G                              (vga_G),                                                              //                        .G
		.vga_B                              (vga_B),                                                              //                        .B
		.vga_pll_ref_clk_clk                (vga_pll_ref_clk_clk),                                                //         vga_pll_ref_clk.clk
		.vga_pll_ref_reset_reset            (vga_pll_ref_reset_reset)                                             //       vga_pll_ref_reset.reset
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.System_PLL_sys_clk_clk                              (system_pll_sys_clk_clk),                                             //                            System_PLL_sys_clk.clk
		.JTAG_UART_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                     //         JTAG_UART_reset_reset_bridge_in_reset.reset
		.Nios2_reset_reset_bridge_in_reset_reset             (rst_controller_001_reset_out_reset),                                 //             Nios2_reset_reset_bridge_in_reset.reset
		.VGA_Subsystem_sys_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                     // VGA_Subsystem_sys_reset_reset_bridge_in_reset.reset
		.Nios2_data_master_address                           (nios2_data_master_address),                                          //                             Nios2_data_master.address
		.Nios2_data_master_waitrequest                       (nios2_data_master_waitrequest),                                      //                                              .waitrequest
		.Nios2_data_master_byteenable                        (nios2_data_master_byteenable),                                       //                                              .byteenable
		.Nios2_data_master_read                              (nios2_data_master_read),                                             //                                              .read
		.Nios2_data_master_readdata                          (nios2_data_master_readdata),                                         //                                              .readdata
		.Nios2_data_master_readdatavalid                     (nios2_data_master_readdatavalid),                                    //                                              .readdatavalid
		.Nios2_data_master_write                             (nios2_data_master_write),                                            //                                              .write
		.Nios2_data_master_writedata                         (nios2_data_master_writedata),                                        //                                              .writedata
		.Nios2_data_master_debugaccess                       (nios2_data_master_debugaccess),                                      //                                              .debugaccess
		.Nios2_instruction_master_address                    (nios2_instruction_master_address),                                   //                      Nios2_instruction_master.address
		.Nios2_instruction_master_waitrequest                (nios2_instruction_master_waitrequest),                               //                                              .waitrequest
		.Nios2_instruction_master_read                       (nios2_instruction_master_read),                                      //                                              .read
		.Nios2_instruction_master_readdata                   (nios2_instruction_master_readdata),                                  //                                              .readdata
		.Nios2_instruction_master_readdatavalid              (nios2_instruction_master_readdatavalid),                             //                                              .readdatavalid
		.VGA_Subsystem_pixel_dma_master_address              (vga_subsystem_pixel_dma_master_address),                             //                VGA_Subsystem_pixel_dma_master.address
		.VGA_Subsystem_pixel_dma_master_waitrequest          (vga_subsystem_pixel_dma_master_waitrequest),                         //                                              .waitrequest
		.VGA_Subsystem_pixel_dma_master_read                 (vga_subsystem_pixel_dma_master_read),                                //                                              .read
		.VGA_Subsystem_pixel_dma_master_readdata             (vga_subsystem_pixel_dma_master_readdata),                            //                                              .readdata
		.VGA_Subsystem_pixel_dma_master_readdatavalid        (vga_subsystem_pixel_dma_master_readdatavalid),                       //                                              .readdatavalid
		.VGA_Subsystem_pixel_dma_master_lock                 (vga_subsystem_pixel_dma_master_lock),                                //                                              .lock
		.Interval_Timer_s1_address                           (mm_interconnect_0_interval_timer_s1_address),                        //                             Interval_Timer_s1.address
		.Interval_Timer_s1_write                             (mm_interconnect_0_interval_timer_s1_write),                          //                                              .write
		.Interval_Timer_s1_readdata                          (mm_interconnect_0_interval_timer_s1_readdata),                       //                                              .readdata
		.Interval_Timer_s1_writedata                         (mm_interconnect_0_interval_timer_s1_writedata),                      //                                              .writedata
		.Interval_Timer_s1_chipselect                        (mm_interconnect_0_interval_timer_s1_chipselect),                     //                                              .chipselect
		.JTAG_UART_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),              //                   JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                //                                              .write
		.JTAG_UART_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                 //                                              .read
		.JTAG_UART_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),             //                                              .readdata
		.JTAG_UART_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),            //                                              .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),          //                                              .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),           //                                              .chipselect
		.Nios2_debug_mem_slave_address                       (mm_interconnect_0_nios2_debug_mem_slave_address),                    //                         Nios2_debug_mem_slave.address
		.Nios2_debug_mem_slave_write                         (mm_interconnect_0_nios2_debug_mem_slave_write),                      //                                              .write
		.Nios2_debug_mem_slave_read                          (mm_interconnect_0_nios2_debug_mem_slave_read),                       //                                              .read
		.Nios2_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_debug_mem_slave_readdata),                   //                                              .readdata
		.Nios2_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_debug_mem_slave_writedata),                  //                                              .writedata
		.Nios2_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_debug_mem_slave_byteenable),                 //                                              .byteenable
		.Nios2_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),                //                                              .waitrequest
		.Nios2_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),                //                                              .debugaccess
		.Pushbuttons_s1_address                              (mm_interconnect_0_pushbuttons_s1_address),                           //                                Pushbuttons_s1.address
		.Pushbuttons_s1_write                                (mm_interconnect_0_pushbuttons_s1_write),                             //                                              .write
		.Pushbuttons_s1_readdata                             (mm_interconnect_0_pushbuttons_s1_readdata),                          //                                              .readdata
		.Pushbuttons_s1_writedata                            (mm_interconnect_0_pushbuttons_s1_writedata),                         //                                              .writedata
		.Pushbuttons_s1_chipselect                           (mm_interconnect_0_pushbuttons_s1_chipselect),                        //                                              .chipselect
		.SD_Card_avalon_sdcard_slave_address                 (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),              //                   SD_Card_avalon_sdcard_slave.address
		.SD_Card_avalon_sdcard_slave_write                   (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),                //                                              .write
		.SD_Card_avalon_sdcard_slave_read                    (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),                 //                                              .read
		.SD_Card_avalon_sdcard_slave_readdata                (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),             //                                              .readdata
		.SD_Card_avalon_sdcard_slave_writedata               (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),            //                                              .writedata
		.SD_Card_avalon_sdcard_slave_byteenable              (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),           //                                              .byteenable
		.SD_Card_avalon_sdcard_slave_waitrequest             (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest),          //                                              .waitrequest
		.SD_Card_avalon_sdcard_slave_chipselect              (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),           //                                              .chipselect
		.SDRAM_s1_address                                    (mm_interconnect_0_sdram_s1_address),                                 //                                      SDRAM_s1.address
		.SDRAM_s1_write                                      (mm_interconnect_0_sdram_s1_write),                                   //                                              .write
		.SDRAM_s1_read                                       (mm_interconnect_0_sdram_s1_read),                                    //                                              .read
		.SDRAM_s1_readdata                                   (mm_interconnect_0_sdram_s1_readdata),                                //                                              .readdata
		.SDRAM_s1_writedata                                  (mm_interconnect_0_sdram_s1_writedata),                               //                                              .writedata
		.SDRAM_s1_byteenable                                 (mm_interconnect_0_sdram_s1_byteenable),                              //                                              .byteenable
		.SDRAM_s1_readdatavalid                              (mm_interconnect_0_sdram_s1_readdatavalid),                           //                                              .readdatavalid
		.SDRAM_s1_waitrequest                                (mm_interconnect_0_sdram_s1_waitrequest),                             //                                              .waitrequest
		.SDRAM_s1_chipselect                                 (mm_interconnect_0_sdram_s1_chipselect),                              //                                              .chipselect
		.SRAM_avalon_sram_slave_address                      (mm_interconnect_0_sram_avalon_sram_slave_address),                   //                        SRAM_avalon_sram_slave.address
		.SRAM_avalon_sram_slave_write                        (mm_interconnect_0_sram_avalon_sram_slave_write),                     //                                              .write
		.SRAM_avalon_sram_slave_read                         (mm_interconnect_0_sram_avalon_sram_slave_read),                      //                                              .read
		.SRAM_avalon_sram_slave_readdata                     (mm_interconnect_0_sram_avalon_sram_slave_readdata),                  //                                              .readdata
		.SRAM_avalon_sram_slave_writedata                    (mm_interconnect_0_sram_avalon_sram_slave_writedata),                 //                                              .writedata
		.SRAM_avalon_sram_slave_byteenable                   (mm_interconnect_0_sram_avalon_sram_slave_byteenable),                //                                              .byteenable
		.SRAM_avalon_sram_slave_readdatavalid                (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid),             //                                              .readdatavalid
		.SysID_control_slave_address                         (mm_interconnect_0_sysid_control_slave_address),                      //                           SysID_control_slave.address
		.SysID_control_slave_readdata                        (mm_interconnect_0_sysid_control_slave_readdata),                     //                                              .readdata
		.VGA_Subsystem_pixel_dma_control_slave_address       (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address),    //         VGA_Subsystem_pixel_dma_control_slave.address
		.VGA_Subsystem_pixel_dma_control_slave_write         (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write),      //                                              .write
		.VGA_Subsystem_pixel_dma_control_slave_read          (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read),       //                                              .read
		.VGA_Subsystem_pixel_dma_control_slave_readdata      (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata),   //                                              .readdata
		.VGA_Subsystem_pixel_dma_control_slave_writedata     (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata),  //                                              .writedata
		.VGA_Subsystem_pixel_dma_control_slave_byteenable    (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable)  //                                              .byteenable
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (system_pll_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (nios2_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (system_pll_reset_source_reset),  // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_debug_reset_request_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),          // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
